// Only for numbers and letters which can be
// displayed well on a seven-segment nixie tube
`define DISP_0 8'b00000011
`define DISP_1 8'b10011111
`define DISP_2 8'b00100101
`define DISP_3 8'b00001101
`define DISP_4 8'b10011001
`define DISP_5 8'b01001001
`define DISP_6 8'b01000001
`define DISP_7 8'b00011111
`define DISP_8 8'b00000001
`define DISP_9 8'b00001001
`define DISP_A 8'b00010001
`define DISP_C 8'b01100011
`define DISP_E 8'b01100001
`define DISP_F 8'b01110001
`define DISP_G 8'b01000011
`define DISP_H 8'b10010001
`define DISP_L 8'b11100001
`define DISP_O 8'b00000011
`define DISP_P 8'b00110001
`define DISP_U 8'b10000011